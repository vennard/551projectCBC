module test();

//some sort of bit swizzzzlers

endmodule:
