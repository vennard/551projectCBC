library verilog;
use verilog.vl_types.all;
entity cbc_dig_tb is
end cbc_dig_tb;
