library verilog;
use verilog.vl_types.all;
entity datapath_control is
end datapath_control;
